`timescale 1ns / 1ps

module CacheInterface(
    input [31:0] ADDR,
    input [31:0] DI,
    input WE,
    output [31:0] DO,
    output RDY
    );


endmodule
